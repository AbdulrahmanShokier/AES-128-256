module round_0 #(parameter BLOCK_LENGTH = 128)
(
    input                         clk,
    input                         rst,  
    input      [BLOCK_LENGTH-1:0] IN,
    input      [BLOCK_LENGTH-1:0] KEY,
    output reg [BLOCK_LENGTH-1:0] OUT,
    output reg           valid
);

wire [127:0] xor_out;

key_add xor_with_k0 (.IN(IN), .KEY(KEY), .OUT(xor_out)); // first step

always@(posedge clk or negedge rst)
begin

    valid <= 1'b0;
    if(!rst)
    begin
        OUT <= 128'b0;
    end

    else
    begin
        OUT <= xor_out;
    end
    
end


always@(negedge clk or negedge rst)
begin
    if(!rst)
    begin
        valid <= 1'b0;
    end

    else
    begin
        valid <= 1'b1;
    end
    
end

endmodule