 module S_box

(
	//Ports declaration.
	
	// Input data to the "Substitute_Bytes" stage statge (1 byte). 
	input      [8-1:0] in_byte,
	
	// Output data from the "Substitute_Bytes" statge (1 byte). 	
	output reg [8-1:0] out_byte
);
  
 //Code starts here
//-----------------------------------------------------------------------------//

  always @ (*)  // Start of the always block.
                // Sensitivity list contains data_in.
  begin
	
		//LUT of "Substitute_Bytes" stage
		case (in_byte) 
		    8'h 00 : out_byte = 8'h 63 ;
			8'h 10 : out_byte = 8'h CA ;
			8'h 20 : out_byte = 8'h B7 ;
			8'h 30 : out_byte = 8'h 04 ;
			8'h 40 : out_byte = 8'h 09 ;
			8'h 50 : out_byte = 8'h 53 ;
			8'h 60 : out_byte = 8'h D0 ;
			8'h 70 : out_byte = 8'h 51 ;
			8'h 80 : out_byte = 8'h CD ;
			8'h 90 : out_byte = 8'h 60 ;
			8'h A0 : out_byte = 8'h E0 ;
			8'h B0 : out_byte = 8'h E7 ;
			8'h C0 : out_byte = 8'h BA ;
			8'h D0 : out_byte = 8'h 70 ;
			8'h E0 : out_byte = 8'h E1 ;
			8'h F0 : out_byte = 8'h 8C ;
			8'h 01 : out_byte = 8'h 7C ;
			8'h 11 : out_byte = 8'h 82 ;
			8'h 21 : out_byte = 8'h FD ;
			8'h 31 : out_byte = 8'h C7 ;
			8'h 41 : out_byte = 8'h 83 ;
			8'h 51 : out_byte = 8'h D1 ;
			8'h 61 : out_byte = 8'h EF ;
			8'h 71 : out_byte = 8'h A3 ;
			8'h 81 : out_byte = 8'h 0C ;
			8'h 91 : out_byte = 8'h 81 ;
			8'h A1 : out_byte = 8'h 32 ;
			8'h B1 : out_byte = 8'h C8 ;
			8'h C1 : out_byte = 8'h 78 ;
			8'h D1 : out_byte = 8'h 3E ;
			8'h E1 : out_byte = 8'h F8 ;
			8'h F1 : out_byte = 8'h A1 ;
			8'h 02 : out_byte = 8'h 77 ;
			8'h 12 : out_byte = 8'h C9 ;
			8'h 22 : out_byte = 8'h 93 ;
			8'h 32 : out_byte = 8'h 23 ;
			8'h 42 : out_byte = 8'h 2C ;
			8'h 52 : out_byte = 8'h 00 ;
			8'h 62 : out_byte = 8'h AA ;
			8'h 72 : out_byte = 8'h 40 ;
			8'h 82 : out_byte = 8'h 13 ;
			8'h 92 : out_byte = 8'h 4F ;
			8'h A2 : out_byte = 8'h 3A ;
			8'h B2 : out_byte = 8'h 37 ;
			8'h C2 : out_byte = 8'h 25 ;
			8'h D2 : out_byte = 8'h B5 ;
			8'h E2 : out_byte = 8'h 98 ;
			8'h F2 : out_byte = 8'h 89 ;
			8'h 03 : out_byte = 8'h 7B ;
			8'h 13 : out_byte = 8'h 7D ;
			8'h 23 : out_byte = 8'h 26 ;
			8'h 33 : out_byte = 8'h C3 ;
			8'h 43 : out_byte = 8'h 1A ;
			8'h 53 : out_byte = 8'h ED ;
			8'h 63 : out_byte = 8'h FB ;
			8'h 73 : out_byte = 8'h 8F ;
			8'h 83 : out_byte = 8'h EC ;
			8'h 93 : out_byte = 8'h DC ;
			8'h A3 : out_byte = 8'h 0A ;
			8'h B3 : out_byte = 8'h 6D ;
			8'h C3 : out_byte = 8'h 2E ;
			8'h D3 : out_byte = 8'h 66 ;
			8'h E3 : out_byte = 8'h 11 ;
			8'h F3 : out_byte = 8'h 0D ;
			8'h 04 : out_byte = 8'h F2 ;
			8'h 14 : out_byte = 8'h FA ;
			8'h 24 : out_byte = 8'h 36 ;
			8'h 34 : out_byte = 8'h 18 ;
			8'h 44 : out_byte = 8'h 1B ;
			8'h 54 : out_byte = 8'h 20 ;
			8'h 64 : out_byte = 8'h 43 ;
			8'h 74 : out_byte = 8'h 92 ;
			8'h 84 : out_byte = 8'h 5F ;
			8'h 94 : out_byte = 8'h 22 ;
			8'h A4 : out_byte = 8'h 49 ;
			8'h B4 : out_byte = 8'h 8D ;
			8'h C4 : out_byte = 8'h 1C ;
			8'h D4 : out_byte = 8'h 48 ;
			8'h E4 : out_byte = 8'h 69 ;
			8'h F4 : out_byte = 8'h BF ;
			8'h 05 : out_byte = 8'h 6B ;
			8'h 15 : out_byte = 8'h 59 ;
			8'h 25 : out_byte = 8'h 3F ;
			8'h 35 : out_byte = 8'h 96 ;
			8'h 45 : out_byte = 8'h 6E ;
			8'h 55 : out_byte = 8'h FC ;
			8'h 65 : out_byte = 8'h 4D ;
			8'h 75 : out_byte = 8'h 9D ;
			8'h 85 : out_byte = 8'h 97 ;
			8'h 95 : out_byte = 8'h 2A ;
			8'h A5 : out_byte = 8'h 06 ;
			8'h B5 : out_byte = 8'h D5 ;
			8'h C5 : out_byte = 8'h A6 ;
			8'h D5 : out_byte = 8'h 03 ;
			8'h E5 : out_byte = 8'h D9 ;
			8'h F5 : out_byte = 8'h E6 ;
			8'h 06 : out_byte = 8'h 6F ;
			8'h 16 : out_byte = 8'h 47 ;
			8'h 26 : out_byte = 8'h F7 ;
			8'h 36 : out_byte = 8'h 05 ;
			8'h 46 : out_byte = 8'h 5A ;
			8'h 56 : out_byte = 8'h B1 ;
			8'h 66 : out_byte = 8'h 33 ;
			8'h 76 : out_byte = 8'h 38 ;
			8'h 86 : out_byte = 8'h 44 ;
			8'h 96 : out_byte = 8'h 90 ;
			8'h A6 : out_byte = 8'h 24 ;
			8'h B6 : out_byte = 8'h 4E ;
			8'h C6 : out_byte = 8'h B4 ;
			8'h D6 : out_byte = 8'h F6 ;
			8'h E6 : out_byte = 8'h 8E ;
			8'h F6 : out_byte = 8'h 42 ;
			8'h 07 : out_byte = 8'h C5 ;
			8'h 17 : out_byte = 8'h F0 ;
			8'h 27 : out_byte = 8'h CC ;
			8'h 37 : out_byte = 8'h 9A ;
			8'h 47 : out_byte = 8'h A0 ;
			8'h 57 : out_byte = 8'h 5B ;
			8'h 67 : out_byte = 8'h 85 ;
			8'h 77 : out_byte = 8'h F5 ;
			8'h 87 : out_byte = 8'h 17 ;
			8'h 97 : out_byte = 8'h 88 ;
			8'h A7 : out_byte = 8'h 5C ;
			8'h B7 : out_byte = 8'h A9 ;
			8'h C7 : out_byte = 8'h C6 ;
			8'h D7 : out_byte = 8'h 0E ;
			8'h E7 : out_byte = 8'h 94 ;
			8'h F7 : out_byte = 8'h 68 ;
			8'h 08 : out_byte = 8'h 30 ;
			8'h 18 : out_byte = 8'h AD ;
			8'h 28 : out_byte = 8'h 34 ;
			8'h 38 : out_byte = 8'h 07 ;
			8'h 48 : out_byte = 8'h 52 ;
			8'h 58 : out_byte = 8'h 6A ;
			8'h 68 : out_byte = 8'h 45 ;
			8'h 78 : out_byte = 8'h BC ;
			8'h 88 : out_byte = 8'h C4 ;
			8'h 98 : out_byte = 8'h 46 ;
			8'h A8 : out_byte = 8'h C2 ;
			8'h B8 : out_byte = 8'h 6C ;
			8'h C8 : out_byte = 8'h E8 ;
			8'h D8 : out_byte = 8'h 61 ;
			8'h E8 : out_byte = 8'h 9B ;
			8'h F8 : out_byte = 8'h 41 ;
			8'h 09 : out_byte = 8'h 01 ;
			8'h 19 : out_byte = 8'h D4 ;
			8'h 29 : out_byte = 8'h A5 ;
			8'h 39 : out_byte = 8'h 12 ;
			8'h 49 : out_byte = 8'h 3B ;
			8'h 59 : out_byte = 8'h CB ;
			8'h 69 : out_byte = 8'h F9 ;
			8'h 79 : out_byte = 8'h B6 ;
			8'h 89 : out_byte = 8'h A7 ;
			8'h 99 : out_byte = 8'h EE ;
			8'h A9 : out_byte = 8'h D3 ;
			8'h B9 : out_byte = 8'h 56 ;
			8'h C9 : out_byte = 8'h DD ;
			8'h D9 : out_byte = 8'h 35 ;
			8'h E9 : out_byte = 8'h 1E ;
			8'h F9 : out_byte = 8'h 99 ;
			8'h 0A : out_byte = 8'h 67 ;
			8'h 1A : out_byte = 8'h A2 ;
			8'h 2A : out_byte = 8'h E5 ;
			8'h 3A : out_byte = 8'h 80 ;
			8'h 4A : out_byte = 8'h D6 ;
			8'h 5A : out_byte = 8'h BE ;
			8'h 6A : out_byte = 8'h 02 ;
			8'h 7A : out_byte = 8'h DA ;
			8'h 8A : out_byte = 8'h 7E ;
			8'h 9A : out_byte = 8'h B8 ;
			8'h AA : out_byte = 8'h AC ;
			8'h BA : out_byte = 8'h F4 ;
			8'h CA : out_byte = 8'h 74 ;
			8'h DA : out_byte = 8'h 57 ;
			8'h EA : out_byte = 8'h 87 ;
			8'h FA : out_byte = 8'h 2D ;
			8'h 0B : out_byte = 8'h 2B ;
			8'h 1B : out_byte = 8'h AF ;
			8'h 2B : out_byte = 8'h F1 ;
			8'h 3B : out_byte = 8'h E2 ;
			8'h 4B : out_byte = 8'h B3 ;
			8'h 5B : out_byte = 8'h 39 ;
			8'h 6B : out_byte = 8'h 7F ;
			8'h 7B : out_byte = 8'h 21 ;
			8'h 8B : out_byte = 8'h 3D ;
			8'h 9B : out_byte = 8'h 14 ;
			8'h AB : out_byte = 8'h 62 ;
			8'h BB : out_byte = 8'h EA ;
			8'h CB : out_byte = 8'h 1F ;
			8'h DB : out_byte = 8'h B9 ;
			8'h EB : out_byte = 8'h E9 ;
			8'h FB : out_byte = 8'h 0F ;
			8'h 0C : out_byte = 8'h FE ;
			8'h 1C : out_byte = 8'h 9C ;
			8'h 2C : out_byte = 8'h 71 ;
			8'h 3C : out_byte = 8'h EB ;
			8'h 4C : out_byte = 8'h 29 ;
			8'h 5C : out_byte = 8'h 4A ;
			8'h 6C : out_byte = 8'h 50 ;
			8'h 7C : out_byte = 8'h 10 ;
			8'h 8C : out_byte = 8'h 64 ;
			8'h 9C : out_byte = 8'h DE ;
			8'h AC : out_byte = 8'h 91 ;
			8'h BC : out_byte = 8'h 65 ;
			8'h CC : out_byte = 8'h 4B ;
			8'h DC : out_byte = 8'h 86 ;
			8'h EC : out_byte = 8'h CE ;
			8'h FC : out_byte = 8'h B0 ;
			8'h 0D : out_byte = 8'h D7 ;
			8'h 1D : out_byte = 8'h A4 ;
			8'h 2D : out_byte = 8'h D8 ;
			8'h 3D : out_byte = 8'h 27 ;
			8'h 4D : out_byte = 8'h E3 ;
			8'h 5D : out_byte = 8'h 4C ;
			8'h 6D : out_byte = 8'h 3C ;
			8'h 7D : out_byte = 8'h FF ;
			8'h 8D : out_byte = 8'h 5D ;
			8'h 9D : out_byte = 8'h 5E ;
			8'h AD : out_byte = 8'h 95 ;
			8'h BD : out_byte = 8'h 7A ;
			8'h CD : out_byte = 8'h BD ;
			8'h DD : out_byte = 8'h C1 ;
			8'h ED : out_byte = 8'h 55 ;
			8'h FD : out_byte = 8'h 54 ;
			8'h 0E : out_byte = 8'h AB ;
			8'h 1E : out_byte = 8'h 72 ;
			8'h 2E : out_byte = 8'h 31 ;
			8'h 3E : out_byte = 8'h B2 ;
			8'h 4E : out_byte = 8'h 2F ;
			8'h 5E : out_byte = 8'h 58 ;
			8'h 6E : out_byte = 8'h 9F ;
			8'h 7E : out_byte = 8'h F3 ;
			8'h 8E : out_byte = 8'h 19 ;
			8'h 9E : out_byte = 8'h 0B ;
			8'h AE : out_byte = 8'h E4 ;
			8'h BE : out_byte = 8'h AE ;
			8'h CE : out_byte = 8'h 8B ;
			8'h DE : out_byte = 8'h 1D ;
			8'h EE : out_byte = 8'h 28 ;
			8'h FE : out_byte = 8'h BB ;
			8'h 0F : out_byte = 8'h 76 ;
			8'h 1F : out_byte = 8'h C0 ;
			8'h 2F : out_byte = 8'h 15 ;
			8'h 3F : out_byte = 8'h 75 ;
			8'h 4F : out_byte = 8'h 84 ;
			8'h 5F : out_byte = 8'h CF ;
			8'h 6F : out_byte = 8'h A8 ;
			8'h 7F : out_byte = 8'h D2 ;
			8'h 8F : out_byte = 8'h 73 ;
			8'h 9F : out_byte = 8'h DB ;
			8'h AF : out_byte = 8'h 79 ;
			8'h BF : out_byte = 8'h 08 ;
			8'h CF : out_byte = 8'h 8A ;
			8'h DF : out_byte = 8'h 9E ;
			8'h EF : out_byte = 8'h DF ;
			8'h FF : out_byte = 8'h 16; 
		endcase // End of case.

end // End of always.
 //-----------------------------------------------------------------------------// 
 
endmodule // End of module.