module gf_multiplier #(
    parameter m = 8
)(
    input              clk,
    input              rst_n,
    input  [m-1 : 0]   op_a,
    input  [m-1 : 0]   op_b,
    output reg [m-1 : 0] result
);

// ═══════════════════════════════════════════════════════════
// LOG TABLE: Maps field element to its logarithm (power of α)
// log_rom[α^i] = i
// log_rom[0] = 0 (undefined, but set to 0 for handling)
// ═══════════════════════════════════════════════════════════
reg [m-1 : 0] log_rom [0:255];

// ═══════════════════════════════════════════════════════════
// EXP TABLE (ANTILOG): Maps power of α to field element
// exp_rom[i] = α^i
// Extended to 510 to avoid modulo operation in lookup
// ═══════════════════════════════════════════════════════════
reg [m-1 : 0] exp_rom [0:510];

// Pipeline registers
reg [m-1 : 0] log_a; 
reg [m-1 : 0] log_b;
reg [m-1 : 0] log_sum;

// Zero detection pipeline
reg zero_a_stage1, zero_b_stage1;
reg zero_result_stage2;
reg zero_result_stage3;

// ═══════════════════════════════════════════════════════════
// ROM INITIALIZATION
// ═══════════════════════════════════════════════════════════
initial begin
    integer i;
    
    // Initialize LOG ROM
    // log_rom[0] = 0 (special case, 0 has no logarithm)
    log_rom[0] = 8'd0;
    log_rom[1] = 8'd0;    // α^0 = 1
    log_rom[2] = 8'd1;    // α^1 = 2
    log_rom[4] = 8'd2;    // α^2 = 4
    log_rom[8] = 8'd3;    // α^3 = 8
    log_rom[16] = 8'd4;   // α^4 = 16
    log_rom[32] = 8'd5;   // α^5 = 32
    log_rom[64] = 8'd6;   // α^6 = 64
    log_rom[128] = 8'd7;  // α^7 = 128
    log_rom[29] = 8'd8;   // α^8 = 29 (reduced by primitive poly)
    log_rom[58] = 8'd9;   // α^9 = 58
    log_rom[116] = 8'd10; // α^10 = 116
    log_rom[232] = 8'd11; // α^11 = 232
    log_rom[205] = 8'd12; // α^12 = 205
    log_rom[135] = 8'd13; // α^13 = 135
    log_rom[19] = 8'd14;  // α^14 = 19
    log_rom[38] = 8'd15;  // α^15 = 38
    log_rom[76] = 8'd16;  // α^16 = 76
    log_rom[152] = 8'd17; // α^17 = 152
    log_rom[45] = 8'd18;  // α^18 = 45
    log_rom[90] = 8'd19;  // α^19 = 90
    log_rom[180] = 8'd20; // α^20 = 180
    log_rom[117] = 8'd21; // α^21 = 117
    log_rom[234] = 8'd22; // α^22 = 234
    log_rom[201] = 8'd23; // α^23 = 201
    log_rom[143] = 8'd24; // α^24 = 143
    log_rom[3] = 8'd25;   // α^25 = 3
    log_rom[6] = 8'd26;   // α^26 = 6
    log_rom[12] = 8'd27;  // α^27 = 12
    log_rom[24] = 8'd28;  // α^28 = 24
    log_rom[48] = 8'd29;  // α^29 = 48
    log_rom[96] = 8'd30;  // α^30 = 96
    log_rom[192] = 8'd31; // α^31 = 192
    log_rom[157] = 8'd32; // α^32 = 157
    log_rom[39] = 8'd33;  // α^33 = 39
    log_rom[78] = 8'd34;  // α^34 = 78
    log_rom[156] = 8'd35; // α^35 = 156
    log_rom[37] = 8'd36;  // α^36 = 37
    log_rom[74] = 8'd37;  // α^37 = 74
    log_rom[148] = 8'd38; // α^38 = 148
    log_rom[53] = 8'd39;  // α^39 = 53
    log_rom[106] = 8'd40; // α^40 = 106
    log_rom[212] = 8'd41; // α^41 = 212
    log_rom[181] = 8'd42; // α^42 = 181
    log_rom[119] = 8'd43; // α^43 = 119
    log_rom[238] = 8'd44; // α^44 = 238
    log_rom[193] = 8'd45; // α^45 = 193
    log_rom[159] = 8'd46; // α^46 = 159
    log_rom[35] = 8'd47;  // α^47 = 35
    log_rom[70] = 8'd48;  // α^48 = 70
    log_rom[140] = 8'd49; // α^49 = 140
    log_rom[5] = 8'd50;   // α^50 = 5
    log_rom[10] = 8'd51;  // α^51 = 10
    log_rom[20] = 8'd52;  // α^52 = 20
    log_rom[40] = 8'd53;  // α^53 = 40
    log_rom[80] = 8'd54;  // α^54 = 80
    log_rom[160] = 8'd55; // α^55 = 160
    log_rom[93] = 8'd56;  // α^56 = 93
    log_rom[186] = 8'd57; // α^57 = 186
    log_rom[105] = 8'd58; // α^58 = 105
    log_rom[210] = 8'd59; // α^59 = 210
    log_rom[185] = 8'd60; // α^60 = 185
    log_rom[111] = 8'd61; // α^61 = 111
    log_rom[222] = 8'd62; // α^62 = 222
    log_rom[161] = 8'd63; // α^63 = 161
    log_rom[95] = 8'd64;  // α^64 = 95
    log_rom[190] = 8'd65; // α^65 = 190
    log_rom[97] = 8'd66;  // α^66 = 97
    log_rom[194] = 8'd67; // α^67 = 194
    log_rom[153] = 8'd68; // α^68 = 153
    log_rom[47] = 8'd69;  // α^69 = 47
    log_rom[94] = 8'd70;  // α^70 = 94
    log_rom[188] = 8'd71; // α^71 = 188
    log_rom[101] = 8'd72; // α^72 = 101
    log_rom[202] = 8'd73; // α^73 = 202
    log_rom[137] = 8'd74; // α^74 = 137
    log_rom[15] = 8'd75;  // α^75 = 15
    log_rom[30] = 8'd76;  // α^76 = 30
    log_rom[60] = 8'd77;  // α^77 = 60
    log_rom[120] = 8'd78; // α^78 = 120
    log_rom[240] = 8'd79; // α^79 = 240
    log_rom[253] = 8'd80; // α^80 = 253
    log_rom[231] = 8'd81; // α^81 = 231
    log_rom[211] = 8'd82; // α^82 = 211
    log_rom[187] = 8'd83; // α^83 = 187
    log_rom[107] = 8'd84; // α^84 = 107
    log_rom[214] = 8'd85; // α^85 = 214
    log_rom[177] = 8'd86; // α^86 = 177
    log_rom[127] = 8'd87; // α^87 = 127
    log_rom[254] = 8'd88; // α^88 = 254
    log_rom[225] = 8'd89; // α^89 = 225
    log_rom[223] = 8'd90; // α^90 = 223
    log_rom[163] = 8'd91; // α^91 = 163
    log_rom[91] = 8'd92;  // α^92 = 91
    log_rom[182] = 8'd93; // α^93 = 182
    log_rom[113] = 8'd94; // α^94 = 113
    log_rom[226] = 8'd95; // α^95 = 226
    log_rom[217] = 8'd96; // α^96 = 217
    log_rom[175] = 8'd97; // α^97 = 175
    log_rom[67] = 8'd98;  // α^98 = 67
    log_rom[134] = 8'd99; // α^99 = 134
    log_rom[17] = 8'd100; // α^100 = 17
    log_rom[34] = 8'd101; // α^101 = 34
    log_rom[68] = 8'd102; // α^102 = 68
    log_rom[136] = 8'd103; // α^103 = 136
    log_rom[13] = 8'd104;  // α^104 = 13
    log_rom[26] = 8'd105;  // α^105 = 26
    log_rom[52] = 8'd106;  // α^106 = 52
    log_rom[104] = 8'd107; // α^107 = 104
    log_rom[208] = 8'd108; // α^108 = 208
    log_rom[189] = 8'd109; // α^109 = 189
    log_rom[103] = 8'd110; // α^110 = 103
    log_rom[206] = 8'd111; // α^111 = 206
    log_rom[129] = 8'd112; // α^112 = 129
    log_rom[31] = 8'd113;  // α^113 = 31
    log_rom[62] = 8'd114;  // α^114 = 62
    log_rom[124] = 8'd115; // α^115 = 124
    log_rom[248] = 8'd116; // α^116 = 248
    log_rom[237] = 8'd117; // α^117 = 237
    log_rom[199] = 8'd118; // α^118 = 199
    log_rom[147] = 8'd119; // α^119 = 147
    log_rom[59] = 8'd120;  // α^120 = 59
    log_rom[118] = 8'd121; // α^121 = 118
    log_rom[236] = 8'd122; // α^122 = 236
    log_rom[197] = 8'd123; // α^123 = 197
    log_rom[151] = 8'd124; // α^124 = 151
    log_rom[51] = 8'd125;  // α^125 = 51
    log_rom[102] = 8'd126; // α^126 = 102
    log_rom[204] = 8'd127; // α^127 = 204
    log_rom[133] = 8'd128; // α^128 = 133
    log_rom[23] = 8'd129;  // α^129 = 23
    log_rom[46] = 8'd130;  // α^130 = 46
    log_rom[92] = 8'd131;  // α^131 = 92
    log_rom[184] = 8'd132; // α^132 = 184
    log_rom[109] = 8'd133; // α^133 = 109
    log_rom[218] = 8'd134; // α^134 = 218
    log_rom[169] = 8'd135; // α^135 = 169
    log_rom[79] = 8'd136;  // α^136 = 79
    log_rom[158] = 8'd137; // α^137 = 158
    log_rom[33] = 8'd138;  // α^138 = 33
    log_rom[66] = 8'd139;  // α^139 = 66
    log_rom[132] = 8'd140; // α^140 = 132
    log_rom[21] = 8'd141;  // α^141 = 21
    log_rom[42] = 8'd142;  // α^142 = 42
    log_rom[84] = 8'd143;  // α^143 = 84
    log_rom[168] = 8'd144; // α^144 = 168
    log_rom[77] = 8'd145;  // α^145 = 77
    log_rom[154] = 8'd146; // α^146 = 154
    log_rom[41] = 8'd147;  // α^147 = 41
    log_rom[82] = 8'd148;  // α^148 = 82
    log_rom[164] = 8'd149; // α^149 = 164
    log_rom[85] = 8'd150;  // α^150 = 85
    log_rom[170] = 8'd151; // α^151 = 170
    log_rom[73] = 8'd152;  // α^152 = 73
    log_rom[146] = 8'd153; // α^153 = 146
    log_rom[57] = 8'd154;  // α^154 = 57
    log_rom[114] = 8'd155; // α^155 = 114
    log_rom[228] = 8'd156; // α^156 = 228
    log_rom[213] = 8'd157; // α^157 = 213
    log_rom[183] = 8'd158; // α^158 = 183
    log_rom[115] = 8'd159; // α^159 = 115
    log_rom[230] = 8'd160; // α^160 = 230
    log_rom[209] = 8'd161; // α^161 = 209
    log_rom[191] = 8'd162; // α^162 = 191
    log_rom[99] = 8'd163;  // α^163 = 99
    log_rom[198] = 8'd164; // α^164 = 198
    log_rom[145] = 8'd165; // α^165 = 145
    log_rom[63] = 8'd166;  // α^166 = 63
    log_rom[126] = 8'd167; // α^167 = 126
    log_rom[252] = 8'd168; // α^168 = 252
    log_rom[229] = 8'd169; // α^169 = 229
    log_rom[215] = 8'd170; // α^170 = 215
    log_rom[179] = 8'd171; // α^171 = 179
    log_rom[123] = 8'd172; // α^172 = 123
    log_rom[246] = 8'd173; // α^173 = 246
    log_rom[241] = 8'd174; // α^174 = 241
    log_rom[255] = 8'd175; // α^175 = 255
    log_rom[227] = 8'd176; // α^176 = 227
    log_rom[219] = 8'd177; // α^177 = 219
    log_rom[171] = 8'd178; // α^178 = 171
    log_rom[75] = 8'd179;  // α^179 = 75
    log_rom[150] = 8'd180; // α^180 = 150
    log_rom[49] = 8'd181;  // α^181 = 49
    log_rom[98] = 8'd182;  // α^182 = 98
    log_rom[196] = 8'd183; // α^183 = 196
    log_rom[149] = 8'd184; // α^184 = 149
    log_rom[55] = 8'd185;  // α^185 = 55
    log_rom[110] = 8'd186; // α^186 = 110
    log_rom[220] = 8'd187; // α^187 = 220
    log_rom[165] = 8'd188; // α^188 = 165
    log_rom[87] = 8'd189;  // α^189 = 87
    log_rom[174] = 8'd190; // α^190 = 174
    log_rom[65] = 8'd191;  // α^191 = 65
    log_rom[130] = 8'd192; // α^192 = 130
    log_rom[25] = 8'd193;  // α^193 = 25
    log_rom[50] = 8'd194;  // α^194 = 50
    log_rom[100] = 8'd195; // α^195 = 100
    log_rom[200] = 8'd196; // α^196 = 200
    log_rom[141] = 8'd197; // α^197 = 141
    log_rom[7] = 8'd198;   // α^198 = 7
    log_rom[14] = 8'd199;  // α^199 = 14
    log_rom[28] = 8'd200;  // α^200 = 28
    log_rom[56] = 8'd201;  // α^201 = 56
    log_rom[112] = 8'd202; // α^202 = 112
    log_rom[224] = 8'd203; // α^203 = 224
    log_rom[221] = 8'd204; // α^204 = 221
    log_rom[167] = 8'd205; // α^205 = 167
    log_rom[83] = 8'd206;  // α^206 = 83
    log_rom[166] = 8'd207; // α^207 = 166
    log_rom[81] = 8'd208;  // α^208 = 81
    log_rom[162] = 8'd209; // α^209 = 162
    log_rom[89] = 8'd210;  // α^210 = 89
    log_rom[178] = 8'd211; // α^211 = 178
    log_rom[121] = 8'd212; // α^212 = 121
    log_rom[242] = 8'd213; // α^213 = 242
    log_rom[249] = 8'd214; // α^214 = 249
    log_rom[239] = 8'd215; // α^215 = 239
    log_rom[195] = 8'd216; // α^216 = 195
    log_rom[155] = 8'd217; // α^217 = 155
    log_rom[43] = 8'd218;  // α^218 = 43
    log_rom[86] = 8'd219;  // α^219 = 86
    log_rom[172] = 8'd220; // α^220 = 172
    log_rom[69] = 8'd221;  // α^221 = 69
    log_rom[138] = 8'd222; // α^222 = 138
    log_rom[9] = 8'd223;   // α^223 = 9
    log_rom[18] = 8'd224;  // α^224 = 18
    log_rom[36] = 8'd225;  // α^225 = 36
    log_rom[72] = 8'd226;  // α^226 = 72
    log_rom[144] = 8'd227; // α^227 = 144
    log_rom[61] = 8'd228;  // α^228 = 61
    log_rom[122] = 8'd229; // α^229 = 122
    log_rom[244] = 8'd230; // α^230 = 244
    log_rom[245] = 8'd231; // α^231 = 245
    log_rom[247] = 8'd232; // α^232 = 247
    log_rom[243] = 8'd233; // α^233 = 243
    log_rom[251] = 8'd234; // α^234 = 251
    log_rom[235] = 8'd235; // α^235 = 235
    log_rom[203] = 8'd236; // α^236 = 203
    log_rom[139] = 8'd237; // α^237 = 139
    log_rom[11] = 8'd238;  // α^238 = 11
    log_rom[22] = 8'd239;  // α^239 = 22
    log_rom[44] = 8'd240;  // α^240 = 44
    log_rom[88] = 8'd241;  // α^241 = 88
    log_rom[176] = 8'd242; // α^242 = 176
    log_rom[125] = 8'd243; // α^243 = 125
    log_rom[250] = 8'd244; // α^244 = 250
    log_rom[233] = 8'd245; // α^245 = 233
    log_rom[207] = 8'd246; // α^246 = 207
    log_rom[131] = 8'd247; // α^247 = 131
    log_rom[27] = 8'd248;  // α^248 = 27
    log_rom[54] = 8'd249;  // α^249 = 54
    log_rom[108] = 8'd250; // α^250 = 108
    log_rom[216] = 8'd251; // α^251 = 216
    log_rom[173] = 8'd252; // α^252 = 173
    log_rom[71] = 8'd253;  // α^253 = 71
    log_rom[142] = 8'd254; // α^254 = 142
    // α^255 = α^0 = 1 (wraps around)

    // Initialize EXP ROM (extended to 510 to avoid modulo)
    exp_rom[0] = 8'd1;    // α^0
    exp_rom[1] = 8'd2;    // α^1
    exp_rom[2] = 8'd4;    // α^2
    exp_rom[3] = 8'd8;    // α^3
    exp_rom[4] = 8'd16;   // α^4
    exp_rom[5] = 8'd32;   // α^5
    exp_rom[6] = 8'd64;   // α^6
    exp_rom[7] = 8'd128;  // α^7
    exp_rom[8] = 8'd29;   // α^8
    exp_rom[9] = 8'd58;   // α^9
    exp_rom[10] = 8'd116; // α^10
    exp_rom[11] = 8'd232; // α^11
    exp_rom[12] = 8'd205; // α^12
    exp_rom[13] = 8'd135; // α^13
    exp_rom[14] = 8'd19;  // α^14
    exp_rom[15] = 8'd38;  // α^15
    exp_rom[16] = 8'd76;  // α^16
    exp_rom[17] = 8'd152; // α^17
    exp_rom[18] = 8'd45;  // α^18
    exp_rom[19] = 8'd90;  // α^19
    exp_rom[20] = 8'd180; // α^20
    exp_rom[21] = 8'd117; // α^21
    exp_rom[22] = 8'd234; // α^22
    exp_rom[23] = 8'd201; // α^23
    exp_rom[24] = 8'd143; // α^24
    exp_rom[25] = 8'd3;   // α^25
    exp_rom[26] = 8'd6;   // α^26
    exp_rom[27] = 8'd12;  // α^27
    exp_rom[28] = 8'd24;  // α^28
    exp_rom[29] = 8'd48;  // α^29
    exp_rom[30] = 8'd96;  // α^30
    exp_rom[31] = 8'd192; // α^31
    exp_rom[32] = 8'd157; // α^32
    exp_rom[33] = 8'd39;  // α^33
    exp_rom[34] = 8'd78;  // α^34
    exp_rom[35] = 8'd156; // α^35
    exp_rom[36] = 8'd37;  // α^36
    exp_rom[37] = 8'd74;  // α^37
    exp_rom[38] = 8'd148; // α^38
    exp_rom[39] = 8'd53;  // α^39
    exp_rom[40] = 8'd106; // α^40
    exp_rom[41] = 8'd212; // α^41
    exp_rom[42] = 8'd181; // α^42
    exp_rom[43] = 8'd119; // α^43
    exp_rom[44] = 8'd238; // α^44
    exp_rom[45] = 8'd193; // α^45
    exp_rom[46] = 8'd159; // α^46
    exp_rom[47] = 8'd35;  // α^47
    exp_rom[48] = 8'd70;  // α^48
    exp_rom[49] = 8'd140; // α^49
    exp_rom[50] = 8'd5;   // α^50
    exp_rom[51] = 8'd10;  // α^51
    exp_rom[52] = 8'd20;  // α^52
    exp_rom[53] = 8'd40;  // α^53
    exp_rom[54] = 8'd80;  // α^54
    exp_rom[55] = 8'd160; // α^55
    exp_rom[56] = 8'd93;  // α^56
    exp_rom[57] = 8'd186; // α^57
    exp_rom[58] = 8'd105; // α^58
    exp_rom[59] = 8'd210; // α^59
    exp_rom[60] = 8'd185; // α^60
    exp_rom[61] = 8'd111; // α^61
    exp_rom[62] = 8'd222; // α^62
    exp_rom[63] = 8'd161; // α^63
    exp_rom[64] = 8'd95;  // α^64
    exp_rom[65] = 8'd190; // α^65
    exp_rom[66] = 8'd97;  // α^66
    exp_rom[67] = 8'd194; // α^67
    exp_rom[68] = 8'd153; // α^68
    exp_rom[69] = 8'd47;  // α^69
    exp_rom[70] = 8'd94;  // α^70
    exp_rom[71] = 8'd188; // α^71
    exp_rom[72] = 8'd101; // α^72
    exp_rom[73] = 8'd202; // α^73
    exp_rom[74] = 8'd137; // α^74
    exp_rom[75] = 8'd15;  // α^75
    exp_rom[76] = 8'd30;  // α^76
    exp_rom[77] = 8'd60;  // α^77
    exp_rom[78] = 8'd120; // α^78
    exp_rom[79] = 8'd240; // α^79
    exp_rom[80] = 8'd253; // α^80
    exp_rom[81] = 8'd231; // α^81
    exp_rom[82] = 8'd211; // α^82
    exp_rom[83] = 8'd187; // α^83
    exp_rom[84] = 8'd107; // α^84
    exp_rom[85] = 8'd214; // α^85
    exp_rom[86] = 8'd177; // α^86
    exp_rom[87] = 8'd127; // α^87
    exp_rom[88] = 8'd254; // α^88
    exp_rom[89] = 8'd225; // α^89
    exp_rom[90] = 8'd223; // α^90
    exp_rom[91] = 8'd163; // α^91
    exp_rom[92] = 8'd91;  // α^92
    exp_rom[93] = 8'd182; // α^93
    exp_rom[94] = 8'd113; // α^94
    exp_rom[95] = 8'd226; // α^95
    exp_rom[96] = 8'd217; // α^96
    exp_rom[97] = 8'd175; // α^97
    exp_rom[98] = 8'd67;  // α^98
    exp_rom[99] = 8'd134; // α^99
    exp_rom[100] = 8'd17;  // α^100
    exp_rom[101] = 8'd34;  // α^101
    exp_rom[102] = 8'd68;  // α^102
    exp_rom[103] = 8'd136; // α^103
    exp_rom[104] = 8'd13;  // α^104
    exp_rom[105] = 8'd26;  // α^105
    exp_rom[106] = 8'd52;  // α^106
    exp_rom[107] = 8'd104; // α^107
    exp_rom[108] = 8'd208; // α^108
    exp_rom[109] = 8'd189; // α^109
    exp_rom[110] = 8'd103; // α^110
    exp_rom[111] = 8'd206; // α^111
    exp_rom[112] = 8'd129; // α^112
    exp_rom[113] = 8'd31;  // α^113
    exp_rom[114] = 8'd62;  // α^114
    exp_rom[115] = 8'd124; // α^115
    exp_rom[116] = 8'd248; // α^116
    exp_rom[117] = 8'd237; // α^117
    exp_rom[118] = 8'd199; // α^118
    exp_rom[119] = 8'd147; // α^119
    exp_rom[120] = 8'd59;  // α^120
    exp_rom[121] = 8'd118; // α^121
    exp_rom[122] = 8'd236; // α^122
    exp_rom[123] = 8'd197; // α^123
    exp_rom[124] = 8'd151; // α^124
    exp_rom[125] = 8'd51;  // α^125
    exp_rom[126] = 8'd102; // α^126
    exp_rom[127] = 8'd204; // α^127
    exp_rom[128] = 8'd133; // α^128
    exp_rom[129] = 8'd23;  // α^129
    exp_rom[130] = 8'd46;  // α^130
    exp_rom[131] = 8'd92;  // α^131
    exp_rom[132] = 8'd184; // α^132
    exp_rom[133] = 8'd109; // α^133
    exp_rom[134] = 8'd218; // α^134
    exp_rom[135] = 8'd169; // α^135
    exp_rom[136] = 8'd79;  // α^136
    exp_rom[137] = 8'd158; // α^137
    exp_rom[138] = 8'd33;  // α^138
    exp_rom[139] = 8'd66;  // α^139
    exp_rom[140] = 8'd132; // α^140
    exp_rom[141] = 8'd21;  // α^141
    exp_rom[142] = 8'd42;  // α^142
    exp_rom[143] = 8'd84;  // α^143
    exp_rom[144] = 8'd168; // α^144
    exp_rom[145] = 8'd77;  // α^145
    exp_rom[146] = 8'd154; // α^146
    exp_rom[147] = 8'd41;  // α^147
    exp_rom[148] = 8'd82;  // α^148
    exp_rom[149] = 8'd164; // α^149
    exp_rom[150] = 8'd85;  // α^150
    exp_rom[151] = 8'd170; // α^151
    exp_rom[152] = 8'd73;  // α^152
    exp_rom[153] = 8'd146; // α^153
    exp_rom[154] = 8'd57;  // α^154
    exp_rom[155] = 8'd114; // α^155
    exp_rom[156] = 8'd228; // α^156
    exp_rom[157] = 8'd213; // α^157
    exp_rom[158] = 8'd183; // α^158
    exp_rom[159] = 8'd115; // α^159
    exp_rom[160] = 8'd230; // α^160
    exp_rom[161] = 8'd209; // α^161
    exp_rom[162] = 8'd191; // α^162
    exp_rom[163] = 8'd99;  // α^163
    exp_rom[164] = 8'd198; // α^164
    exp_rom[165] = 8'd145; // α^165
    exp_rom[166] = 8'd63;  // α^166
    exp_rom[167] = 8'd126; // α^167
    exp_rom[168] = 8'd252; // α^168
    exp_rom[169] = 8'd229; // α^169
    exp_rom[170] = 8'd215; // α^170
    exp_rom[171] = 8'd179; // α^171
    exp_rom[172] = 8'd123; // α^172
    exp_rom[173] = 8'd246; // α^173
    exp_rom[174] = 8'd241; // α^174
    exp_rom[175] = 8'd255; // α^175
    exp_rom[176] = 8'd227; // α^176
    exp_rom[177] = 8'd219; // α^177
    exp_rom[178] = 8'd171; // α^178
    exp_rom[179] = 8'd75;  // α^179
    exp_rom[180] = 8'd150; // α^180
    exp_rom[181] = 8'd49;  // α^181
    exp_rom[182] = 8'd98;  // α^182
    exp_rom[183] = 8'd196; // α^183
    exp_rom[184] = 8'd149; // α^184
    exp_rom[185] = 8'd55;  // α^185
    exp_rom[186] = 8'd110; // α^186
    exp_rom[187] = 8'd220; // α^187
    exp_rom[188] = 8'd165; // α^188
    exp_rom[189] = 8'd87;  // α^189
    exp_rom[190] = 8'd174; // α^190
    exp_rom[191] = 8'd65;  // α^191
    exp_rom[192] = 8'd130; // α^192
    exp_rom[193] = 8'd25;  // α^193
    exp_rom[194] = 8'd50;  // α^194
    exp_rom[195] = 8'd100; // α^195
    exp_rom[196] = 8'd200; // α^196
    exp_rom[197] = 8'd141; // α^197
    exp_rom[198] = 8'd7;   // α^198
    exp_rom[199] = 8'd14;  // α^199
    exp_rom[200] = 8'd28;  // α^200
    exp_rom[201] = 8'd56;  // α^201
    exp_rom[202] = 8'd112; // α^202
    exp_rom[203] = 8'd224; // α^203
    exp_rom[204] = 8'd221; // α^204
    exp_rom[205] = 8'd167; // α^205
    exp_rom[206] = 8'd83;  // α^206
    exp_rom[207] = 8'd166; // α^207
    exp_rom[208] = 8'd81;  // α^208
    exp_rom[209] = 8'd162; // α^209
    exp_rom[210] = 8'd89;  // α^210
    exp_rom[211] = 8'd178; // α^211
    exp_rom[212] = 8'd121; // α^212
    exp_rom[213] = 8'd242; // α^213
    exp_rom[214] = 8'd249; // α^214
    exp_rom[215] = 8'd239; // α^215
    exp_rom[216] = 8'd195; // α^216
    exp_rom[217] = 8'd155; // α^217
    exp_rom[218] = 8'd43;  // α^218
    exp_rom[219] = 8'd86;  // α^219
    exp_rom[220] = 8'd172; // α^220
    exp_rom[221] = 8'd69;  // α^221
    exp_rom[222] = 8'd138; // α^222
    exp_rom[223] = 8'd9;   // α^223
    exp_rom[224] = 8'd18;  // α^224
    exp_rom[225] = 8'd36;  // α^225
    exp_rom[226] = 8'd72;  // α^226
    exp_rom[227] = 8'd144; // α^227
    exp_rom[228] = 8'd61;  // α^228
    exp_rom[229] = 8'd122; // α^229
    exp_rom[230] = 8'd244; // α^230
    exp_rom[231] = 8'd245; // α^231
    exp_rom[232] = 8'd247; // α^232
    exp_rom[233] = 8'd243; // α^233
    exp_rom[234] = 8'd251; // α^234
    exp_rom[235] = 8'd235; // α^235
    exp_rom[236] = 8'd203; // α^236
    exp_rom[237] = 8'd139; // α^237
    exp_rom[238] = 8'd11;  // α^238
    exp_rom[239] = 8'd22;  // α^239
    exp_rom[240] = 8'd44;  // α^240
    exp_rom[241] = 8'd88;  // α^241
    exp_rom[242] = 8'd176; // α^242
    exp_rom[243] = 8'd125; // α^243
    exp_rom[244] = 8'd250; // α^244
    exp_rom[245] = 8'd233; // α^245
    exp_rom[246] = 8'd207; // α^246
    exp_rom[247] = 8'd131; // α^247
    exp_rom[248] = 8'd27;  // α^248
    exp_rom[249] = 8'd54;  // α^249
    exp_rom[250] = 8'd108; // α^250
    exp_rom[251] = 8'd216; // α^251
    exp_rom[252] = 8'd173; // α^252
    exp_rom[253] = 8'd71;  // α^253
    exp_rom[254] = 8'd142; // α^254
    
    // Duplicate entries for extended table (255-510)
    // This avoids modulo operation: exp_rom[i+255] = exp_rom[i]
    for (i = 255; i < 511; i = i + 1) begin
        exp_rom[i] = exp_rom[i - 255];
    end
end

// ═══════════════════════════════════════════════════════════
// PIPELINE STAGES
// ═══════════════════════════════════════════════════════════
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        log_a <= 8'd0;
        log_b <= 8'd0;
        log_sum <= 8'd0;
        result <= 8'd0;
        
        zero_a_stage1 <= 1'b0;
        zero_b_stage1 <= 1'b0;
        zero_result_stage2 <= 1'b0;
        zero_result_stage3 <= 1'b0;
    end
    else begin
        // Stage 1: Log table lookup + zero detection
        log_a <= log_rom[op_a];
        log_b <= log_rom[op_b];
        zero_a_stage1 <= (op_a == 8'd0);
        zero_b_stage1 <= (op_b == 8'd0);
        
        // Stage 2: Add logarithms
        log_sum <= log_a + log_b;
        zero_result_stage2 <= zero_a_stage1 | zero_b_stage1;
        
        // Stage 3: Antilog lookup + zero handling
        zero_result_stage3 <= zero_result_stage2;
        if (zero_result_stage2)
            result <= 8'd0;  // If either operand was 0, result is 0
        else
            result <= exp_rom[log_sum];  // Normal case
    end
end

endmodule