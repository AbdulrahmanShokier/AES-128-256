`timescale 1us/1us 

module Key_Gen_TB(); 

/////////////////////////////////////////////////
/////////////////// Parameters //////////////////
/////////////////////////////////////////////////

parameter KEY_LENGTH = 128; 
parameter CLK_PER = 10; 


/////////////////////////////////////////////////
///////////////// Test values ///////////////////
/////////////////////////////////////////////////

reg [KEY_LENGTH-1:0] MainKey = 128'h2B7E151628AED2A6ABF7158809CF4F3C;
reg [KEY_LENGTH-1:0] LastSubKey = 128'hD014F9A8C9EE2589E13F0CC8B6630CA6;


/////////////////////////////////////////////////
//////////////// DUT Signals ////////////////////
/////////////////////////////////////////////////

 reg 					RST_tb; 
 reg 					CLK_tb; 
 reg  [KEY_LENGTH-1:0] 	M_KEY_tb; 		
 reg 					En_tb; 		
 wire [KEY_LENGTH-1:0] 	subKey_curr_tb; 

 
/////////////////////////////////////////////////
//////////////// Initial block //////////////////
/////////////////////////////////////////////////

initial
begin 
	
	RST_tb = 1'b1; 
	CLK_tb = 1'b0;
	M_KEY_tb = MainKey; 
	
	#CLK_PER; 
	RST_tb = 1'b0; 
	#CLK_PER; 
	RST_tb = 1'b1;
	
	#(2*CLK_PER);
	En_tb = 1'b1; 
	
	#(10*CLK_PER);		// only 10 as k0 is output with RST not the clock edge  	
	En_tb = 1'b0; 
	
	if(subKey_curr_tb == LastSubKey)
		$display("PASSED!"); 
	
	#(5*CLK_PER); 
	$stop; 
end 




/////////////////////////////////////////////////
/////////////////// Tasks ///////////////////////
/////////////////////////////////////////////////




/////////////////////////////////////////////////
///////////////// Clock Generator ///////////////
/////////////////////////////////////////////////

always #(CLK_PER/2) CLK_tb = ~CLK_tb; 


/////////////////////////////////////////////////
////////////// DUT Instantiations ///////////////
/////////////////////////////////////////////////

Key_Gen DUT(
.RST(RST_tb), 
.CLK(CLK_tb), 
.M_KEY(M_KEY_tb), 		
.En(En_tb), 		
.subKey_curr(subKey_curr_tb)
); 



endmodule 